000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000777777770000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000022220000000000000000000
000000000000000007700700000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000111100000000000000000000000
000000000000000000250200000000000000000000000000000000000111100000000000
000007007001111000000000012210000000000001221000000000000000000000000000
000000000000000000000000000000011110000000000000000000000000000000000000
000001111000000000000000000000000000011110000000000000000000000000000111
000000000000000000000000000440400000444400000000000000000002200000000006
111111111111111111111111111111111111111111111111111111111111111111111111
